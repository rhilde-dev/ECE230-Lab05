module top(
  input [6:0] sw,
  output [1:0] led
)
  //TODO: feed inputs into circuitA
  //TODO: feed inputs into circuitB
  //find out how to add wires

endmodule
