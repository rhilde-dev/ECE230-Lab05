module top(
  input [6:0] sw,
  output [1:0] led
)

  wire w1;
  
  //TODO: feed inputs into circuit
  //TODO: feed inputs into circuitB
  //find out how to add wires

endmodule
